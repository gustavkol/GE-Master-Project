package tta0_params is
end tta0_params;
