package tta0_params is
  constant fu_lsu_dataw : integer := 32;
  constant fu_lsu_addrw : integer := 8;
end tta0_params;
