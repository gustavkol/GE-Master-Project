library IEEE;
use IEEE.Std_Logic_1164.all;
use std.textio.all;
use ieee.numeric_std.all;

entity testbench is
end testbench;

architecture behav of testbench is

  --  Declaration and binding of the component that will be instantiated.
   component fu_under_test
      port(
      t1data    : in std_logic_vector(31 downto 0);
      t1load    : in  std_logic;
      t2data    : in std_logic_vector(31 downto 0);
      t2load    : in  std_logic;
      r1data    : out std_logic_vector(31 downto 0);
      t1opcode  : in std_logic_vector(2 downto 0);
      glock     : in  std_logic;
      rstx      : in  std_logic;
      clk       : in  std_logic);
   end component;


   for tested_fu_0 : fu_under_test use entity work.fu_algo;

  --  Specify registers for the ports.
   signal t1data        : std_logic_vector(31 downto 0);
   signal t1load        : std_logic_vector(1-1 downto 0);
   signal t2data        : std_logic_vector(31 downto 0);
   signal t2load        : std_logic_vector(1-1 downto 0);
   signal r1data        : std_logic_vector(31 downto 0);
   signal t1opcode      : std_logic_vector(2 downto 0);
   signal glock : std_logic;
   signal rstx  : std_logic;
   signal clk   : std_logic;


begin
  --  Map ports of the FU to registers.
   tested_fu_0  :       fu_under_test
      port map (
         t1data => t1data,
         t1load => t1load(0),
         t2data => t2data,
         t2load => t2load(0),
         r1data => r1data,
         t1opcode => t1opcode,
         clk => clk,
         rstx => rstx,
         glock => glock);
  process

    -- Arrays for stimulus.
      type t1data_data_array is array (natural range <>) of
         std_logic_vector(31 downto 0);

      constant t1data_data : t1data_data_array :=
      ("00000000000000000001001110001000",       -- @0 = 5000 (compare_and_iter_f)
       "00000000000000000001001110001000",       -- @1 = 5000 (compare_and_iter_f)
       "00000000000000000011101010011000",       -- @2 = 15000 (compare_and_iter_f)
       "00000000000000000011101010011000",       -- @3 = 15000 (compare_and_iter_f)
       "00000000000000000110000110101000",       -- @4 = 25000 (compare_and_iter_f)
       "11111111111111111110110001111000",       -- @5 = -5000 (compare_and_iter_f)
       "11111111111111111110110001111000",       -- @6 = -5000 (compare_and_iter_f)
       "11111111111111111100010101101000",       -- @7 = -15000 (compare_and_iter_f)
       "11111111111111111100010101101000",       -- @8 = -15000 (compare_and_iter_f)
       "11111111111111111001111001011000",       -- @9 = -25000 (compare_and_iter_f)
       "00000000000000000010111011100000",       -- @10 = 12 000 (compare_and_iter_int)
       "00000000000000000000000000000000",
       "00000000000000000100111000100000",       -- @11 = 20 000 (compare_and_iter_int)
       "00000000000000000000000000000000",
       "00000000000000000111010100110000",       -- @12 = 30 000 (compare_and_iter_int)
       "00000000000000000000000000000000",
       "00000000000000001010010000010000",       -- @13 = 42 000 (compare_and_iter_int)
       "00000000000000000000000000000000",
       "00000000000000001110101001100000",       -- @14 = 60 000 (compare_and_iter_int)
       "00000000000000000000000000000000",
       "00000000000000011110100001001000",       -- @15 = 125 000 (compare_and_iter_int)
       "00000000000000000000000000000000",
       "00000000000000101011111100100000",       -- @16 = 180 000 (compare_and_iter_int)
       "00000000000000000000000000000000",
       "00000000000000110101101101100000",       -- @17 = 220 000 (compare_and_iter_int)
       "00000000000000000000000000000000",
       "11111111111111111011000111100000",       -- @18 = -20 000 (compare_and_iter_int)
       "00000000000000000000000000000000",
       "11111111111111110001010110100000",       -- @19 = -60 000 (compare_and_iter_int)
       "00000000000000000000000000000000",
       "00001000010101001011101101001110",       -- @20 = 139770702
       "00101111110000000001101000011111",       -- @21 = 801118751
       "10011010100011001011111101001000",       -- @22 = 2592915272
       "01100000010011010111100001011111",       -- @23 = 1615689823
       "00001110001111011100100011011000",       -- @24 = 238930136
       "11111110010001101111100010110101",       -- @25 = 4266064053
       "11110100010110110100110010000011",       -- @26 = 4099624067
       "11111000110011100011111001101000",       -- @27 = 4174265960
       "10010110111011001000001011111000",       -- @28 = 2532082424
       "10011100111000000001100010011110",       -- @29 = 2631932062
       "11100110101000100101110010000111",       -- @30 = 3869400199
       "01000001010011001111101010101011",       -- @31 = 1095563947
       "11000010011000100011100011110111",       -- @32 = 3261217015
       "01100101111111111001011110011110",       -- @33 = 1711249310
       "01101011000100101000010101010000",       -- @34 = 1796375888
       "01011100101011011011000001001001",       -- @35 = 1554886729
       "00010101101110000011001010001011",       -- @36 = 364393099
       "11001011100011100001010111101111",       -- @37 = 3415086575
       "11101111000110010111100100011011",       -- @38 = 4011424027
       "10011000010010011110110001111111",       -- @39 = 2554981503
       "01110111100100011101000011011111",       -- @40 = 2006044895
       "00111110011111111111110000000010",       -- @41 = 1048574978
       "01101011110111100001011000101010",       -- @42 = 1809716778
       "10010000111011110001000101100000",       -- @43 = 2431586656
       "00101101010111110010110001000010",       -- @44 = 761211970
       "10100110110000010101101001111010",       -- @45 = 2797689466
       "11000111100011000101110011111111",       -- @46 = 3347864831
       "00100100110010110110001100101110",       -- @47 = 617308974
       "11101110101100101111101001010000",       -- @48 = 4004706896
       "00011000100011001011110110001001",       -- @49 = 411876745
       "01110010011001001111010101001100",       -- @50 = 1919219020
       "10011101001010000011111010010011",       -- @51 = 2636660371
       "00001100111110001110111101000101",       -- @52 = 217640773
       "01001011010101001011001011000111",       -- @53 = 1263841991
       "11011000111110001101100001111010",       -- @54 = 3640187002
       "00010111010010001010110011000110",       -- @55 = 390638790
       "11100110000000101011100000110001",       -- @56 = 3858937905
       "10100110000011011001001000010101",       -- @57 = 2785907221
       "11110010111011011111100110010111",       -- @58 = 4075682199
       "01011001000000111010001011101010",       -- @59 = 1493410538
       "00001000000101001111111001100101",       -- @60 = 135593573
       "01110110011001111000110010000111",       -- @61 = 1986497671
       "11110101111101111010001010100101",       -- @62 = 4126646949
       "10000000111010011000100010111111",       -- @63 = 2162788543
       "10011000001111100000100110100100",       -- @64 = 2554202532
       "10011010000111011101000010101000",       -- @65 = 2585645224
       "10110111100101011110011010110101",       -- @66 = 3080054453
       "01001001001000000100001101000001",       -- @67 = 1226851137
       "01000001100000110100000110111001",       -- @68 = 1099121081
       "01101110100000010010010000000011",       -- @69 = 1853957123
       "01010101010100001111110111100011",       -- @70 = 1431371235
       "10011000000011000111001001110111",       -- @71 = 2550952567
       "01011111100011001011011111110110",       -- @72 = 1603057654
       "00011000001011110110001110110001",       -- @73 = 405758897
       "01100101010000000001001010010111",       -- @74 = 1698697879
       "01101101011000000101111001110010",       -- @75 = 1835032178
       "11111110010011011101010011110110",       -- @76 = 4266513654
       "10101101010000010000100010100001",       -- @77 = 2906720417
       "11101010100001010000101111100111",       -- @78 = 3934587879
       "00100100001011101001110110010101",       -- @79 = 607034773
       "00000000000000000000000000000000");      -- @80 = 0

      type t2data_data_array is array (natural range <>) of
         std_logic_vector(31 downto 0);

      constant t2data_data : t2data_data_array :=
      ("00000000010011100010000000010000",       -- @0 = 5120016 (compare_and_iter_f)
       "00000000010011100010000000011000",       -- @1 = 5120024 (compare_and_iter_f)
       "00000000010011100010000000010000",       -- @2 = 5120016 (compare_and_iter_f)
       "00000000010011100010000000011000",       -- @3 = 5120024 (compare_and_iter_f)
       "00000000010011100010000000011000",       -- @4 = 5120024 (compare_and_iter_f)
       "00000000010011100010000000010000",       -- @5 = 5120016 (compare_and_iter_f)
       "00000000010011100010000000011000",       -- @6 = 5120024 (compare_and_iter_f)
       "00000000010011100010000000010000",       -- @7 = 5120016 (compare_and_iter_f)
       "00000000010011100010000000011000",       -- @8 = 5120024 (compare_and_iter_f)
       "00000000010011100010000000011000",       -- @9 = 5120024 (compare_and_iter_f)
       "00000000000000000110000110101000",       -- @10 = 25000 (compare_and_iter_int)
       "00000000000000000000000000000000",
       "00000000000000000110000110101000",       -- @11 = 25000 (compare_and_iter_int)
       "00000000000000000000000000000000",
       "00000000000000000110000110101000",       -- @12 = 25000 (compare_and_iter_int)
       "00000000000000000000000000000000",
       "00000000000000000110000110101000",       -- @13 = 25000 (compare_and_iter_int)
       "00000000000000000000000000000000",
       "00000000000000000110000110101000",       -- @14 = 25000 (compare_and_iter_int)
       "00000000000000000000000000000000",
       "00000000000000000110000110101000",       -- @15 = 25000 (compare_and_iter_int)
       "00000000000000000000000000000000",
       "00000000000000000110000110101000",       -- @16 = 25000 (compare_and_iter_int)
       "00000000000000000000000000000000",
       "00000000000000000110000110101000",       -- @17 = 25000 (compare_and_iter_int)
       "00000000000000000000000000000000",
       "00000000000000000110000110101000",       -- @18 = 25000 (compare_and_iter_int)
       "00000000000000000000000000000000",
       "00000000000000000110000110101000",       -- @19 = 25000 (compare_and_iter_int)
       "00000000000000000000000000000000",
       "01111101010001100001110000110001",       -- @20 = 2101746737
       "01100010000100001010000110000011",       -- @21 = 1645257091
       "11111110101010100011110010111100",       -- @22 = 4272569532
       "01110110010100011001100100010110",       -- @23 = 1985059094
       "10000101000110100000110010101110",       -- @24 = 2233076910
       "11001011011000001100101001111101",       -- @25 = 3412118141
       "01000001101011101010000110000110",       -- @26 = 1101963654
       "11110111111011011111100011100001",       -- @27 = 4159568097
       "01000000011100111011010001001101",       -- @28 = 1081324621
       "11101110110000000000010110001011",       -- @29 = 4005561739
       "10100101011101001100110110101011",       -- @30 = 2775895467
       "10100110001111001101001011011110",       -- @31 = 2789003998
       "00001000001111010011111000110011",       -- @32 = 138231347
       "00001010000011110101101001001001",       -- @33 = 168778313
       "00010011100111011010111010110111",       -- @34 = 329100983
       "01001110000110011111111001000111",       -- @35 = 1310326343
       "10111000000100100101101010011010",       -- @36 = 3088210586
       "10011110110100101000101001101111",       -- @37 = 2664598127
       "10111011011100101111001000010101",       -- @38 = 3144872469
       "10001001101000010111000010001010",       -- @39 = 2309058698
       "10011010011110000101110110111111",       -- @40 = 2591579583
       "01111110110011101011101000110010",       -- @41 = 2127477298
       "01100010001011001000000010000100",       -- @42 = 1647083652
       "10011001011110110000001000100000",       -- @43 = 2574975520
       "00100110000011010110111101011101",       -- @44 = 638414685
       "11100010110100010101011000011110",       -- @45 = 3805369886
       "01110111001001000010111100110111",       -- @46 = 1998860087
       "00001000000010001000111000010010",       -- @47 = 134778386
       "11010011111110100100110001101001",       -- @48 = 3556396137
       "00110110001101101101101110000010",       -- @49 = 909564802
       "10000000111110011100000011110000",       -- @50 = 2163851504
       "00100001110100101101110000011000",       -- @51 = 567467032
       "10101110111100011001111100101000",       -- @52 = 2935070504
       "01001100100100011111111110011000",       -- @53 = 1284636568
       "11010100110101111110110110001100",       -- @54 = 3570920844
       "01110010100110011110101111101100",       -- @55 = 1922690028
       "11100011101111101011011011011010",       -- @56 = 3820926682
       "10010111101101110100001000011001",       -- @57 = 2545369625
       "10101010011000011011101010010001",       -- @58 = 2858531473
       "01001011001101001100001000111111",       -- @59 = 1261748799
       "01011011000011101000011100110000",       -- @60 = 1527678768
       "10000001110000101010111010100111",       -- @61 = 2177019559
       "11101110000110010100110010011000",       -- @62 = 3994635416
       "11100101101001001010101110110010",       -- @63 = 3852774322
       "00111011111001100010100010000011",       -- @64 = 1004939395
       "10001000101001100111101110000110",       -- @65 = 2292611974
       "01111110001101010011011110001000",       -- @66 = 2117416840
       "11110110000100011001111101000100",       -- @67 = 4128350020
       "00101100110101100010101001110000",       -- @68 = 752233072
       "11011000000010100010001010111001",       -- @69 = 3624542905
       "11101000101100010010010001110010",       -- @70 = 3903923314
       "10100000101011110000100101111001",       -- @71 = 2695825785
       "00000000010110100100001001010001",       -- @72 = 5915217
       "00110110101101100100110111100001",       -- @73 = 917917153
       "00011111000011001010110001111111",       -- @74 = 520924287
       "10110111110111010000100110110011",       -- @75 = 3084716467
       "00111000100110110000010110100110",       -- @76 = 949683622
       "11110111110011101110110000010011",       -- @77 = 4157533203
       "00001100010000001001010110110011",       -- @78 = 205559219
       "11111100011101101001000111110000",       -- @79 = 4235629040
       "00000000000000000000000000000000");      -- @80 = 0


    -- Opcodes for each clock cycle.
      type t1opcode_data_array is array (natural range <>) of
         std_logic_vector(2 downto 0);

      constant t1opcode_data : t1opcode_data_array :=
      ("001",    -- @0 = 1 (compare_and_iter_f)
       "001",    -- @1 = 1 (compare_and_iter_f)
       "001",    -- @2 = 1 (compare_and_iter_f)
       "001",    -- @3 = 1 (compare_and_iter_f)
       "001",    -- @4 = 1 (compare_and_iter_f)
       "001",    -- @5 = 1 (compare_and_iter_f)
       "001",    -- @6 = 1 (compare_and_iter_f)
       "001",    -- @7 = 1 (compare_and_iter_f)
       "001",    -- @8 = 1 (compare_and_iter_f)
       "001",    -- @9 = 1 (compare_and_iter_f)

       "010",    -- @10 = 2 (compare_and_iter_int)
       "000",
       "010",    -- @11 = 2 (compare_and_iter_int)
       "000",
       "010",    -- @12 = 2 (compare_and_iter_int)
       "000",
       "010",    -- @13 = 2 (compare_and_iter_int)
       "000",
       "010",    -- @14 = 2 (compare_and_iter_int)
       "000",
       "010",    -- @15 = 2 (compare_and_iter_int)
       "000",
       "010",    -- @16 = 2 (compare_and_iter_int)
       "000",
       "010",    -- @17 = 2 (compare_and_iter_int)
       "000",
       "010",    -- @18 = 2 (compare_and_iter_int)
       "000",
       "010",    -- @19 = 2 (compare_and_iter_int)
       "000",

       "100",    -- @20 = 4 (mask_add)
       "100",    -- @21 = 4 (mask_add)
       "100",    -- @22 = 4 (mask_add)
       "100",    -- @23 = 4 (mask_add)
       "100",    -- @24 = 4 (mask_add)
       "100",    -- @25 = 4 (mask_add)
       "100",    -- @26 = 4 (mask_add)
       "100",    -- @27 = 4 (mask_add)
       "100",    -- @28 = 4 (mask_add)
       "100",    -- @29 = 4 (mask_add)
       "101",    -- @30 = 5 (shift_add)
       "101",    -- @31 = 5 (shift_add)
       "101",    -- @32 = 5 (shift_add)
       "101",    -- @33 = 5 (shift_add)
       "101",    -- @34 = 5 (shift_add)
       "101",    -- @35 = 5 (shift_add)
       "101",    -- @36 = 5 (shift_add)
       "101",    -- @37 = 5 (shift_add)
       "101",    -- @38 = 5 (shift_add)
       "101",    -- @39 = 5 (shift_add)
       "000",    -- @40 = 0 (add)
       "000",    -- @41 = 0 (add)
       "000",    -- @42 = 0 (add)
       "000",    -- @43 = 0 (add)
       "000",    -- @44 = 0 (add)
       "000",    -- @45 = 0 (add)
       "000",    -- @46 = 0 (add)
       "000",    -- @47 = 0 (add)
       "000",    -- @48 = 0 (add)
       "000",    -- @49 = 0 (add)
       "110",    -- @50 = 6 (shift_sub)
       "110",    -- @51 = 6 (shift_sub)
       "110",    -- @52 = 6 (shift_sub)
       "110",    -- @53 = 6 (shift_sub)
       "110",    -- @54 = 6 (shift_sub)
       "110",    -- @55 = 6 (shift_sub)
       "110",    -- @56 = 6 (shift_sub)
       "110",    -- @57 = 6 (shift_sub)
       "110",    -- @58 = 6 (shift_sub)
       "110",    -- @59 = 6 (shift_sub)
       "111",    -- @60 = 7 (sub)
       "111",    -- @61 = 7 (sub)
       "111",    -- @62 = 7 (sub)
       "111",    -- @63 = 7 (sub)
       "111",    -- @64 = 7 (sub)
       "111",    -- @65 = 7 (sub)
       "111",    -- @66 = 7 (sub)
       "111",    -- @67 = 7 (sub)
       "111",    -- @68 = 7 (sub)
       "111",    -- @69 = 7 (sub)
       "011",    -- @70 = 3 (inc_comp_next)
       "011",    -- @71 = 3 (inc_comp_next)
       "011",    -- @72 = 3 (inc_comp_next)
       "011",    -- @73 = 3 (inc_comp_next)
       "011",    -- @74 = 3 (inc_comp_next)
       "011",    -- @75 = 3 (inc_comp_next)
       "011",    -- @76 = 3 (inc_comp_next)
       "011",    -- @77 = 3 (inc_comp_next)
       "011",    -- @78 = 3 (inc_comp_next)
       "011",    -- @79 = 3 (inc_comp_next)
       "011");   -- @80 = 3 (inc_comp_next)

    -- Load signals for each cycle
      type t1load_data_array is array (natural range <>) of
         std_logic_vector(0 downto 0);

      constant t1load_data : t1load_data_array :=
      ("1",      -- @0 = 1 (compare_and_iter_f)
       "1",      -- @1 = 1 (compare_and_iter_f)
       "1",      -- @2 = 1 (compare_and_iter_f)
       "1",      -- @3 = 1 (compare_and_iter_f)
       "1",      -- @4 = 1 (compare_and_iter_f)
       "1",      -- @5 = 1 (compare_and_iter_f)
       "1",      -- @6 = 1 (compare_and_iter_f)
       "1",      -- @7 = 1 (compare_and_iter_f)
       "1",      -- @8 = 1 (compare_and_iter_f)
       "1",      -- @9 = 1 (compare_and_iter_f)
       "1",      -- @10 = 1 (compare_and_iter_int)
       "0",
       "1",      -- @11 = 1 (compare_and_iter_int)
       "0",
       "1",      -- @12 = 1 (compare_and_iter_int)
       "0",
       "1",      -- @13 = 1 (compare_and_iter_int)
       "0",
       "1",      -- @14 = 1 (compare_and_iter_int)
       "0",
       "1",      -- @15 = 1 (compare_and_iter_int)
       "0",
       "1",      -- @16 = 1 (compare_and_iter_int)
       "0",
       "1",      -- @17 = 1 (compare_and_iter_int)
       "0",
       "1",      -- @18 = 1 (compare_and_iter_int)
       "0",
       "1",      -- @19 = 1 (compare_and_iter_int)
       "0",
       "1",      -- @20 = 1
       "1",      -- @21 = 1
       "1",      -- @22 = 1
       "1",      -- @23 = 1
       "1",      -- @24 = 1
       "1",      -- @25 = 1
       "1",      -- @26 = 1
       "1",      -- @27 = 1
       "1",      -- @28 = 1
       "1",      -- @29 = 1
       "1",      -- @30 = 1
       "1",      -- @31 = 1
       "1",      -- @32 = 1
       "1",      -- @33 = 1
       "1",      -- @34 = 1
       "1",      -- @35 = 1
       "1",      -- @36 = 1
       "1",      -- @37 = 1
       "1",      -- @38 = 1
       "1",      -- @39 = 1
       "1",      -- @40 = 1
       "1",      -- @41 = 1
       "1",      -- @42 = 1
       "1",      -- @43 = 1
       "1",      -- @44 = 1
       "1",      -- @45 = 1
       "1",      -- @46 = 1
       "1",      -- @47 = 1
       "1",      -- @48 = 1
       "1",      -- @49 = 1
       "1",      -- @50 = 1
       "1",      -- @51 = 1
       "1",      -- @52 = 1
       "1",      -- @53 = 1
       "1",      -- @54 = 1
       "1",      -- @55 = 1
       "1",      -- @56 = 1
       "1",      -- @57 = 1
       "1",      -- @58 = 1
       "1",      -- @59 = 1
       "1",      -- @60 = 1
       "1",      -- @61 = 1
       "1",      -- @62 = 1
       "1",      -- @63 = 1
       "1",      -- @64 = 1
       "1",      -- @65 = 1
       "1",      -- @66 = 1
       "1",      -- @67 = 1
       "1",      -- @68 = 1
       "1",      -- @69 = 1
       "1",      -- @70 = 1
       "1",      -- @71 = 1
       "1",      -- @72 = 1
       "1",      -- @73 = 1
       "1",      -- @74 = 1
       "1",      -- @75 = 1
       "1",      -- @76 = 1
       "1",      -- @77 = 1
       "1",      -- @78 = 1
       "1",      -- @79 = 1
       "0");     -- @80 = 0

      type t2load_data_array is array (natural range <>) of
         std_logic_vector(0 downto 0);

      constant t2load_data : t2load_data_array :=
      ("1",      -- @0 = 1 (compare_and_iter_f)
       "1",      -- @1 = 1 (compare_and_iter_f)
       "1",      -- @2 = 1 (compare_and_iter_f)
       "1",      -- @3 = 1 (compare_and_iter_f)
       "1",      -- @4 = 1 (compare_and_iter_f)
       "1",      -- @5 = 1 (compare_and_iter_f)
       "1",      -- @6 = 1 (compare_and_iter_f)
       "1",      -- @7 = 1 (compare_and_iter_f)
       "1",      -- @8 = 1 (compare_and_iter_f)
       "1",      -- @9 = 1 (compare_and_iter_f)
       "1",      -- @10 = 1 (compare_and_iter_int)
       "0",
       "1",      -- @12 = 1 (compare_and_iter_int)
       "0",
       "1",      -- @14 = 1 (compare_and_iter_int)
       "0",
       "1",      -- @16 = 1 (compare_and_iter_int)
       "0",
       "1",      -- @18 = 1 (compare_and_iter_int)
       "0",
       "1",      -- @20 = 1 (compare_and_iter_int)
       "0",
       "1",      -- @22 = 1 (compare_and_iter_int)
       "0",
       "1",      -- @24 = 1 (compare_and_iter_int)
       "0",
       "1",      -- @26 = 1 (compare_and_iter_int)
       "0",
       "1",      -- @28 = 1 (compare_and_iter_int)
       "0",
       "1",      -- @29 = 1
       "1",      -- @21 = 1
       "1",      -- @22 = 1
       "1",      -- @23 = 1
       "1",      -- @24 = 1
       "1",      -- @25 = 1
       "1",      -- @26 = 1
       "1",      -- @27 = 1
       "1",      -- @28 = 1
       "1",      -- @29 = 1
       "1",      -- @30 = 1
       "1",      -- @31 = 1
       "1",      -- @32 = 1
       "1",      -- @33 = 1
       "1",      -- @34 = 1
       "1",      -- @35 = 1
       "1",      -- @36 = 1
       "1",      -- @37 = 1
       "1",      -- @38 = 1
       "1",      -- @39 = 1
       "1",      -- @40 = 1
       "1",      -- @41 = 1
       "1",      -- @42 = 1
       "1",      -- @43 = 1
       "1",      -- @44 = 1
       "1",      -- @45 = 1
       "1",      -- @46 = 1
       "1",      -- @47 = 1
       "1",      -- @48 = 1
       "1",      -- @49 = 1
       "1",      -- @50 = 1
       "1",      -- @51 = 1
       "1",      -- @52 = 1
       "1",      -- @53 = 1
       "1",      -- @54 = 1
       "1",      -- @55 = 1
       "1",      -- @56 = 1
       "1",      -- @57 = 1
       "1",      -- @58 = 1
       "1",      -- @59 = 1
       "1",      -- @60 = 1
       "1",      -- @61 = 1
       "1",      -- @62 = 1
       "1",      -- @63 = 1
       "1",      -- @64 = 1
       "1",      -- @65 = 1
       "1",      -- @66 = 1
       "1",      -- @67 = 1
       "1",      -- @68 = 1
       "1",      -- @69 = 1
       "1",      -- @70 = 1
       "1",      -- @71 = 1
       "1",      -- @72 = 1
       "1",      -- @73 = 1
       "1",      -- @74 = 1
       "1",      -- @75 = 1
       "1",      -- @76 = 1
       "1",      -- @77 = 1
       "1",      -- @78 = 1
       "1",      -- @79 = 1
       "0");     -- @80 = 0


    -- Arrays for expected outputs for each output port.
      type r1data_data_array is array (natural range <>) of
         std_logic_vector(31 downto 0);

      constant r1data_data : r1data_data_array :=
      ("00000000000000000000000000000000",       -- @0 = 0  
       "00000000000000000000000000010000",       -- @1 = 16 (compare_and_iter_f)
       "00000000000000000000000000011000",       -- @2 = 24 (compare_and_iter_f)
       "00000000001001110010100000010100",       -- @3 = 2566164  (compare_and_iter_f)
       "00000000001001110010110000011100",       -- @4 = 2567196 (compare_and_iter_f)
       "00000000010011100111100000100000",       -- @5 = 5142560 (compare_and_iter_f)
       "00000000000000000000000000010000",       -- @6 = 16 (compare_and_iter_f)
       "00000000000000000000000000011000",       -- @7 = 24 (compare_and_iter_f)
       "11111111110110001111100000001100",       -- @8 = -2557940  (compare_and_iter_f)
       "11111111110110001111010000010100",       -- @9 = -2558956 (compare_and_iter_f)
       "11111111101100100000100000010000",       -- @10 = -5109744    (compare_and_iter_f)
       "11111111101100100000100000010000",       -- @11 = -5109744 (compare_and_iter_f)
       "00000000000000000000000000000000",       -- @12 = 0    (compare_and_iter_int)
       "00000000000000000000000000000000",       
       "00000000001100001101010100000100",       -- @14 = 3200260    (compare_and_iter_int)
       "00000000001100001101010100000100",       
       "00000000011000011010110000001000",       -- @16 = 6401032    (compare_and_iter_int)
       "00000000011000011010110000001000",       
       "00000000100100101000010100001100",       -- @18 = 9602316    (compare_and_iter_int)
       "00000000100100101000010100001100",       
       "00000000110000110110000000010000",       -- @20 = 12804112  (compare_and_iter_int)
       "00000000110000110110000000010000",       
       "00000001101101111100010100100100",       -- @22 = 28820772 (compare_and_iter_int)
       "00000001101101111100010100100100",       
       "00000010101011000101110000111000",       -- @24 = 44850232    (compare_and_iter_int)
       "00000010101011000101110000111000",       
       "00000011001111110011010101000100",       -- @26 = 54474052 (compare_and_iter_int)
       "00000011001111110011010101000100",       
       "11111111110011110010110111111100",       -- @28 = -3199492     (compare_and_iter_int)
       "11111111110011110010110111111100",       
       "11111111001111001100000011110000",       -- @29 = -12795664    (compare_and_iter_int)
       "01111101010001100001110001111111",       -- @21 = 2101746815
       "01100010000100001010000110100010",       -- @22 = 1645257122
       "11111110101010100011110100000100",       -- @23 = 4272569604
       "01110110010100011001100101110101",       -- @24 = 1985059189
       "10000101000110100000110010000110",       -- @25 = 2233076870
       "11001011011000001100101000110010",       -- @26 = 3412118066
       "01000001101011101010000100001001",       -- @27 = 1101963529
       "11110111111011011111100101001001",       -- @28 = 4159568201
       "01000000011100111011010001000101",       -- @29 = 1081324613
       "11101110110000000000010100101001",       -- @30 = 4005561641
       "10100101010110110111000000000111",       -- @31 = 2774233095
       "10100110011111100001111111011000",       -- @32 = 2793283544
       "00000111111111111010000001101011",       -- @33 = 134193259
       "00001010011101010101100111100000",       -- @34 = 175462880
       "00010100000010001100000100111100",       -- @35 = 336118076
       "01001110011101101010101111110111",       -- @36 = 1316400119
       "10111000001010000001001011001100",       -- @37 = 3089633996
       "10011110100111100001100010000100",       -- @38 = 2661161092
       "10111011011000100000101110001110",       -- @39 = 3143764878
       "10001001001110011011101001110110",       -- @40 = 2302261878
       "00010010000010100010111010011110",       -- @41 = 302657182
       "10111101010011101011011000110100",       -- @42 = 3176052276
       "11001110000010101001011010101110",       -- @43 = 3456800430
       "00101010011010100001001110000000",       -- @44 = 711594880
       "01010011011011001001101110011111",       -- @45 = 1399626655
       "10001001100100101011000010011000",       -- @46 = 2308092056
       "00111110101100001000110000110110",       -- @47 = 1051757622
       "00101100110100111111000101000000",       -- @48 = 752087360
       "11000010101011010100011010111001",       -- @49 = 3266135737
       "01001110110000111001100100001011",       -- @50 = 1321441547
       "10000000100001110101101111111011",       -- @51 = 2156354555
       "00100010001101011011001111011010",       -- @52 = 573944794
       "10101110111001001010011000111001",       -- @53 = 2934220345
       "01001100010001101010101011100110",       -- @54 = 1279699686
       "11010100111111101111010010110100",       -- @55 = 3573478580
       "01110010100000101010001101000000",       -- @56 = 1921164096
       "11100011110110001011010000100010",       -- @57 = 3822629922
       "10011000000100010011010010000111",       -- @58 = 2551264391
       "10101010011011101100110010011000",       -- @59 = 2859388056
       "01001010110110111011111010011101",       -- @60 = 1255915165
       "10101101000001100111011100110101",       -- @61 = 2902882101
       "11110100101001001101110111100000",       -- @62 = 4104445408
       "00000111110111100101011000001101",       -- @63 = 132011533
       "10011011010001001101110100001101",       -- @64 = 2604981517
       "01011100010101111110000100100001",       -- @65 = 1549263137
       "00010001011101110101010100100010",       -- @66 = 293033250
       "00111001011000001010111100101101",       -- @67 = 962637613
       "01010011000011101010001111111101",       -- @68 = 1393468413
       "00010100101011010001011101001001",       -- @69 = 346888009
       "10010110011101110000000101001010",       -- @70 = 2524381514
       "10000011111011101011010011111111",       -- @71 = 2213459199
       "01010110101011100101111110000101",       -- @72 = 1454268293
       "01100000010000010011110010011000",       -- @73 = 1614888088
       "10000101100110111111111101110011",       -- @74 = 2241593203
       "10100011010110010110101110010101",       -- @75 = 2740546453
       "11111101101001100100101100001100",       -- @76 = 4255533836
       "01101111100000111110000001000010",       -- @77 = 1870913602
       "10111101101000110011000001111011",       -- @78 = 3181588603
       "00000011000001100011011101001101",       -- @79 = 50739021
       "00101011010000010111100110110101");      -- @80 = 725711285

      constant IGNORE_OUTPUT_COUNT : integer := 1;
      constant TOTAL_CYCLE_COUNT : integer := 90;


     variable current_cycle : integer;
  begin

    -- Initialize the clock signal.
    clk <= '0';

    -- Reset active to initialize regs
    rstx <= '0';
    wait for 1 ns;

    -- Release reset.
    rstx <= '1';
    -- Global lock off.
    glock <= '0';


    for current_cycle in 0 to TOTAL_CYCLE_COUNT - 1 loop

    -- The actual test bench code.
      t1data <= t1data_data(current_cycle);
      t1load <= t1load_data(current_cycle);
      t2data <= t2data_data(current_cycle);
      t2load <= t2load_data(current_cycle);
      t1opcode <= t1opcode_data(current_cycle);

      if current_cycle >= IGNORE_OUTPUT_COUNT then
         assert r1data = r1data_data(current_cycle)
            report lf & "TCE Assert: Verification failed at cycle " & integer'image(current_cycle) & " for output 0"
            & " actual: " & integer'image(to_integer(signed(r1data)))
            & " expected: " & integer'image(to_integer(signed(r1data_data(current_cycle))))  severity error;

      end if;

      -- Generate a clock pulse.
      -- TODO: Generate the clock in a separate component.
      wait for 1 ns;
      clk <= not clk;
      wait for 1 ns;
      clk <= not clk;

    end loop;  -- current_cycle

    -- Ends the simulation (at least in case of ghdl).
    wait;
  end process;
end behav;