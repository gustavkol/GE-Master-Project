library IEEE;
use IEEE.Std_Logic_1164.all;
use std.textio.all;
use ieee.numeric_std.all;

entity testbench is
end testbench;

architecture behav of testbench is

  --  Declaration and binding of the component that will be instantiated.
   component fu_under_test
      port(
      t1data    : in std_logic_vector(31 downto 0);
      t1load    : in  std_logic;
      t2data    : in std_logic_vector(31 downto 0);
      t2load    : in  std_logic;
      r1data    : out std_logic_vector(31 downto 0);
      t1opcode  : in std_logic_vector(2 downto 0);
      glock     : in  std_logic;
      rstx      : in  std_logic;
      clk       : in  std_logic);
   end component;


   for tested_fu_0 : fu_under_test use entity work.fu_algo_frac;

  --  Specify registers for the ports.
   signal t1data        : std_logic_vector(31 downto 0);
   signal t1load        : std_logic_vector(1-1 downto 0);
   signal t2data        : std_logic_vector(31 downto 0);
   signal t2load        : std_logic_vector(1-1 downto 0);
   signal r1data        : std_logic_vector(31 downto 0);
   signal t1opcode      : std_logic_vector(2 downto 0);
   signal glock : std_logic;
   signal rstx  : std_logic;
   signal clk   : std_logic;


begin
  --  Map ports of the FU to registers.
   tested_fu_0  :       fu_under_test
      port map (
         t1data => t1data,
         t1load => t1load(0),
         t2data => t2data,
         t2load => t2load(0),
         r1data => r1data,
         t1opcode => t1opcode,
         clk => clk,
         rstx => rstx,
         glock => glock);
  process

    -- Arrays for stimulus.
      type t1data_data_array is array (natural range <>) of
         std_logic_vector(31 downto 0);

      constant t1data_data : t1data_data_array :=
      ("00000000000000000001001110001000",       -- @0 = 5000 (compare_and_iter_f)
       "00000000000000000001001110001000",       -- @1 = 5000 (compare_and_iter_f)
       "11111111111111111110110001111000",       -- @2 = -5000 (compare_and_iter_f)
       "00000000000000000011101010011000",       -- @3 = 15000 (compare_and_iter_f)
       "00000000000000000011101010011000",       -- @4 = 15000 (compare_and_iter_f)
       "11111111111111111100010101101000",       -- @5 = -15000 (compare_and_iter_f)
       "00000000000000000110000110101000",       -- @6 = 25000 (compare_and_iter_f)
       "11111111111111111110110001111000",       -- @7 = -5000 (compare_and_iter_f)
       "11111111111111111110110001111000",       -- @8 = -5000 (compare_and_iter_f)
       "11111111111111111100010101101000",       -- @9 = -15000 (compare_and_iter_f)
       "11111111111111111100010101101000",       -- @10 = -15000 (compare_and_iter_f)
       "11111111111111111100010101101000",       -- @11 = -15000 (compare_and_iter_f)
       "00000000000000000011101010011000",       -- @12 = 15000 (compare_and_iter_f)
       "11110000010011110001100010111111",       -- @10 = 4031715519
       "01011110000001000101010111011111",       -- @11 = 1577342431
       "10111011100000110111001011111100",       -- @12 = 3145954044
       "10101011000111101110110001101011",       -- @13 = 2870930539
       "01111011100101101100010000111000",       -- @14 = 2073478200
       "10101000110010101001110001110010",       -- @15 = 2831850610
       "10110010001101000111001111001001",       -- @16 = 2989781961
       "00101111100100010010100011011011",       -- @17 = 798042331
       "10010111000111001000011111111101",       -- @18 = 2535229437
       "01010110000010110001011011100101",       -- @19 = 1443567333
       "00110101110001001011010000000101",       -- @20 = 902083589
       "01111100000011001100001110100101",       -- @21 = 2081211301
       "10010110000101010100000101011110",       -- @22 = 2517975390
       "11010001111001111011100010001011",       -- @23 = 3521624203
       "11000101010010011000111101001010",       -- @24 = 3309932362
       "10010110011010010011110110111100",       -- @25 = 2523479484
       "11101100000000100110111100110000",       -- @26 = 3959582512
       "00000010000110101010000010010000",       -- @27 = 35299472
       "01100010101100110010101111110000",       -- @28 = 1655909360
       "00110001000001000101010110001010",       -- @29 = 822367626
       "10100100100101100110011001000011",       -- @30 = 2761320003
       "01001111010111011000101100111111",       -- @31 = 1331530559
       "01100010010001000101110100010110",       -- @32 = 1648647446
       "01101010000000001100110100001011",       -- @33 = 1778437387
       "10100101011010001000100001001110",       -- @34 = 2775091278
       "11000100101110010001010100101110",       -- @35 = 3300463918
       "10001100111010011101000011010100",       -- @36 = 2364133588
       "00111011110001110001000110101011",       -- @37 = 1002901931
       "11110101110100011101000111101111",       -- @38 = 4124168687
       "10001000100011011100100010011110",       -- @39 = 2290993310
       "11110101010001111000111010001111",       -- @40 = 4115107471
       "11110101100111111000010000011001",       -- @41 = 4120871961
       "00110101100101111111111001111010",       -- @42 = 899153530
       "01010111101110011001001001010100",       -- @43 = 1471779412
       "11110100011010010111000010010001",       -- @44 = 4100550801
       "10011000101101001111011110111000",       -- @45 = 2561996728
       "00110001000110111100111110011011",       -- @46 = 823906203
       "10010100101110011111000001110010",       -- @47 = 2495213682
       "11110100110111000110000010100110",       -- @48 = 4108083366
       "11101000111101111110111111000100",       -- @49 = 3908562884
       "11111111001001100100100111101010",       -- @50 = 4280699370
       "10111001101100010010011110110010",       -- @51 = 3115394994
       "01101000100100101010010010000101",       -- @52 = 1754440837
       "00100000111100001101100110010001",       -- @53 = 552655249
       "11010111101000101000000110000111",       -- @54 = 3617751431
       "01010111100101011001111110011100",       -- @55 = 1469423516
       "11010010110110001001001001010000",       -- @56 = 3537408592
       "01100010000011011101011011010101",       -- @57 = 1645074133
       "11010010000110011011110101100101",       -- @58 = 3524902245
       "01110000010111011101100111011000",       -- @59 = 1885198808
       "01101010010100111101100001000000",       -- @60 = 1783879744
       "10101000101011100111001011101001",       -- @61 = 2830004969
       "11000111110011001110111110001101",       -- @62 = 3352096653
       "10001000011101100100010101010010",       -- @63 = 2289452370
       "10000001011111111101100010101011",       -- @64 = 2172639403
       "10110111001011110000000100100011",       -- @65 = 3073311011
       "10011110111010100001111010111111",       -- @66 = 2666143423
       "01000001100011001011101111110001",       -- @67 = 1099742193
       "11000010011001011011000010101111",       -- @68 = 3261444271
       "01100100101101100011010001101110",       -- @69 = 1689662574
       "00000000000000000000000000000000",       -- @70 = 0 (compare_and_iter_f_init)
       "00000000000000000000000000000100",       -- @71 = 0.25 (compare_and_iter_f_init)
       "00000000000000000000000000010100",       -- @72 = 1.25 (compare_and_iter_f_init)
       "00000000000000000000000000011000",       -- @73 = 1.5 (compare_and_iter_f_init)
       "00000000000000000000000000101000",       -- @74 = 2.5 (compare_and_iter_f_init)
       "00000000000000000000000001001000",       -- @75 = 4.5 (compare_and_iter_f_init)
       "00000000000000000000000001000100",       -- @76 = 4.25 (compare_and_iter_f_init)
       "00000000000000000000000000100000",       -- @77 = 2 (compare_and_iter_f_init)
       "00000000000000000000000001001000",       -- @78 = 4.5 (compare_and_iter_f_init)
       "00000000000000000000000000111100",       -- @79 = 3.75 (compare_and_iter_f_init)
       "00000000000000000000000000000000");      -- @80 = 0

      type t2data_data_array is array (natural range <>) of
         std_logic_vector(31 downto 0);

      constant t2data_data : t2data_data_array :=
      ("00000000010011100010000000010000",       -- @0 = 5120016 (compare_and_iter_f)
       "00000000010011100010000000011000",       -- @1 = 5120024 (compare_and_iter_f)
       "00000000010011100010000011110000",       -- @2 = 5120240 (compare_and_iter_f)
       "00000000010011100010000000010000",       -- @3 = 5120016 (compare_and_iter_f)
       "00000000010011100010000000011000",       -- @4 = 5120024 (compare_and_iter_f)
       "00000000010011100010000011110000",       -- @5 = 5120240 (compare_and_iter_f)
       "00000000010011100010000000100000",       -- @6 = 5120032 (compare_and_iter_f)
       "00000000010011100010000000010000",       -- @7 = 5120016 (compare_and_iter_f)
       "00000000010011100010000000011000",       -- @8 = 5120024 (compare_and_iter_f)
       "00000000010011100010000000010000",       -- @9 = 5120016 (compare_and_iter_f)
       "00000000010011100010000000011000",       -- @10 = 5120024 (compare_and_iter_f)
       "00000000010011100010000000100000",       -- @11 = 5120032 (compare_and_iter_f)
       "00000000010011100010000011101000",       -- @12 = 5120232 (compare_and_iter_f)
       "11010000100111011000110010011110",       -- @13 = 3499986078
       "11000100000111101010010110111111",       -- @11 = 3290342847
       "10111001011111110111101110110111",       -- @12 = 3112139703
       "11000011110100110110101111100010",       -- @13 = 3285412834
       "00101011101010011001110101001001",       -- @14 = 732536137
       "00010110001001001110001011010011",       -- @15 = 371516115
       "11001001010001011100101011000010",       -- @16 = 3376794306
       "10011001000000100101000111101110",       -- @17 = 2567066094
       "11100010101001111010100000001010",       -- @18 = 3802638346
       "01101101101110110011001000110110",       -- @19 = 1840984630
       "00010001100010101001101010001000",       -- @20 = 294296200
       "10010111110100000101110010100110",       -- @21 = 2547014822
       "10001110000110000011000110111111",       -- @22 = 2383950271
       "01101001111001011011111011001100",       -- @23 = 1776664268
       "01110001001011010111001111000111",       -- @24 = 1898804167
       "00011000011101101000111110001010",       -- @25 = 410423178
       "11010011111100100100101011100111",       -- @26 = 3555871463
       "01001001011010001000000100011111",       -- @27 = 1231585567
       "10000011101100110101001000111000",       -- @28 = 2209567288
       "11110110111111101011100100101001",       -- @29 = 4143888681
       "01010000111001000111100010010011",       -- @30 = 1357150355
       "00101110100110111100010001010010",       -- @31 = 781960274
       "01001011111011010000000011011010",       -- @32 = 1273823450
       "11000111010100010111100010000111",       -- @33 = 3344005255
       "11101010110110111010001000100101",       -- @34 = 3940262437
       "01111110011110111110100100100010",       -- @35 = 2122049826
       "11010010011011010011100001000000",       -- @36 = 3530373184
       "11111110011011011101001011010000",       -- @37 = 4268610256
       "10110100011000010010111111111001",       -- @38 = 3026268153
       "11111011000100101000001011101010",       -- @39 = 4212294378
       "01101010000001101101010100101111",       -- @40 = 1778832687
       "10000001111011101100011100111010",       -- @41 = 2179909434
       "00110110010111100000101001100001",       -- @42 = 912132705
       "11110100101001110000010100011011",       -- @43 = 4104586523
       "10100000111001111011010010010010",       -- @44 = 2699539602
       "01001000100000000111001011011111",       -- @45 = 1216377567
       "01011101011100000011001111111010",       -- @46 = 1567634426
       "10111111101001110111000001001110",       -- @47 = 3215421518
       "11001101111001100110010000000000",       -- @48 = 3454428160
       "01110110111000011000101110101011",       -- @49 = 1994492843
       "00001001010001100010011010011000",       -- @50 = 155592344
       "00100111001011011000110111010010",       -- @51 = 657296850
       "11101011000111011101001111111000",       -- @52 = 3944600568
       "00000011111000111001111010010101",       -- @53 = 65248917
       "10000111011000011011010001110000",       -- @54 = 2271327344
       "11010110101001001010101001001100",       -- @55 = 3601115724
       "01001000100110010100001111110010",       -- @56 = 1218003954
       "01110001000101100100101110111111",       -- @57 = 1897286591
       "00011100000111000011110111110101",       -- @58 = 471612917
       "01110010000011001101011100111001",       -- @59 = 1913444153
       "01000000111010010111000100010111",       -- @60 = 1089040663
       "10001101100011101000110001010010",       -- @61 = 2374929490
       "00110101000101100100110000011010",       -- @62 = 890653722
       "10100000111001001111110111011111",       -- @63 = 2699361759
       "00111001110010011111111111110011",       -- @64 = 969539571
       "10011110111100000100000010010100",       -- @65 = 2666545300
       "10011110001110110100010000010011",       -- @66 = 2654684179
       "00101000101101101110000011000101",       -- @67 = 683073733
       "10011100100001001011111100000100",       -- @68 = 2625945348
       "00101110111010101111010100001000",       -- @69 = 787150088
       "00000000000000000000000000010000",       -- @70 = 16 (compare_and_iter_f_init)
       "00000000000000000000000000100100",       -- @71 = 36 (compare_and_iter_f_init)
       "00000000000000000000000000011100",       -- @72 = 28 (compare_and_iter_f_init)
       "11111111111111111111111111010100",       -- @73 = -44 (compare_and_iter_f_init)
       "00000000000000000000000001011000",       -- @74 = 88 (compare_and_iter_f_init)
       "11111111111111111111111111000100",       -- @75 = -60 (compare_and_iter_f_init)
       "00000000000000000000000001000000",       -- @76 = 64 (compare_and_iter_f_init)
       "11111111111111111111111111110000",       -- @77 = -16 (compare_and_iter_f_init)
       "00000000000000000000000001001100",       -- @78 = 76 (compare_and_iter_f_init)
       "00000000000000000000000000100100",       -- @79 = 36 (compare_and_iter_f_init)
       "00000000000000000000000000000000");      -- @80 = 0


    -- Opcodes for each clock cycle.
      type t1opcode_data_array is array (natural range <>) of
         std_logic_vector(2 downto 0);

      constant t1opcode_data : t1opcode_data_array :=
      ("001",    -- @0 = 1 (compare_and_iter_f)
       "001",    -- @1 = 1 (compare_and_iter_f)
       "001",    -- @2 = 1 (compare_and_iter_f)
       "001",    -- @3 = 1 (compare_and_iter_f)
       "001",    -- @4 = 1 (compare_and_iter_f)
       "001",    -- @5 = 1 (compare_and_iter_f)
       "001",    -- @6 = 1 (compare_and_iter_f)
       "001",    -- @7 = 1 (compare_and_iter_f)
       "001",    -- @8 = 1 (compare_and_iter_f)
       "001",    -- @9 = 1 (compare_and_iter_f)
       "001",    -- @10 = 1 (compare_and_iter_f)
       "001",    -- @11 = 1 (compare_and_iter_f)
       "001",    -- @12 = 1 (compare_and_iter_f)
       "011",    -- @10 = 3 (mask_add)
       "011",    -- @11 = 3 (mask_add)
       "011",    -- @12 = 3 (mask_add)
       "011",    -- @13 = 3 (mask_add)
       "011",    -- @14 = 3 (mask_add)
       "011",    -- @15 = 3 (mask_add)
       "011",    -- @16 = 3 (mask_add)
       "011",    -- @17 = 3 (mask_add)
       "011",    -- @18 = 3 (mask_add)
       "011",    -- @19 = 3 (mask_add)
       "101",    -- @20 = 5 (shift_add)
       "101",    -- @21 = 5 (shift_add)
       "101",    -- @22 = 5 (shift_add)
       "101",    -- @23 = 5 (shift_add)
       "101",    -- @24 = 5 (shift_add)
       "101",    -- @25 = 5 (shift_add)
       "101",    -- @26 = 5 (shift_add)
       "101",    -- @27 = 5 (shift_add)
       "101",    -- @28 = 5 (shift_add)
       "101",    -- @29 = 5 (shift_add)
       "000",    -- @30 = 0 (add)
       "000",    -- @31 = 0 (add)
       "000",    -- @32 = 0 (add)
       "000",    -- @33 = 0 (add)
       "000",    -- @34 = 0 (add)
       "000",    -- @35 = 0 (add)
       "000",    -- @36 = 0 (add)
       "000",    -- @37 = 0 (add)
       "000",    -- @38 = 0 (add)
       "000",    -- @39 = 0 (add)
       "110",    -- @40 = 6 (shift_sub)
       "110",    -- @41 = 6 (shift_sub)
       "110",    -- @42 = 6 (shift_sub)
       "110",    -- @43 = 6 (shift_sub)
       "110",    -- @44 = 6 (shift_sub)
       "110",    -- @45 = 6 (shift_sub)
       "110",    -- @46 = 6 (shift_sub)
       "110",    -- @47 = 6 (shift_sub)
       "110",    -- @48 = 6 (shift_sub)
       "110",    -- @49 = 6 (shift_sub)
       "111",    -- @50 = 7 (sub)
       "111",    -- @51 = 7 (sub)
       "111",    -- @52 = 7 (sub)
       "111",    -- @53 = 7 (sub)
       "111",    -- @54 = 7 (sub)
       "111",    -- @55 = 7 (sub)
       "111",    -- @56 = 7 (sub)
       "111",    -- @57 = 7 (sub)
       "111",    -- @58 = 7 (sub)
       "111",    -- @59 = 7 (sub)
       "100",    -- @60 = 4 (merge)
       "100",    -- @61 = 4 (merge)
       "100",    -- @62 = 4 (merge)
       "100",    -- @63 = 4 (merge)
       "100",    -- @64 = 4 (merge)
       "100",    -- @65 = 4 (merge)
       "100",    -- @66 = 4 (merge)
       "100",    -- @67 = 4 (merge)
       "100",    -- @68 = 4 (merge)
       "100",    -- @69 = 4 (merge)
       "010",    -- @70 = 2 (compare_and_iter_f_init)
       "010",    -- @71 = 2 (compare_and_iter_f_init)
       "010",    -- @72 = 2 (compare_and_iter_f_init)
       "010",    -- @73 = 2 (compare_and_iter_f_init)
       "010",    -- @74 = 2 (compare_and_iter_f_init)
       "010",    -- @75 = 2 (compare_and_iter_f_init)
       "010",    -- @76 = 2 (compare_and_iter_f_init)
       "010",    -- @77 = 2 (compare_and_iter_f_init)
       "010",    -- @78 = 2 (compare_and_iter_f_init)
       "010",    -- @79 = 2 (compare_and_iter_f_init)
       "010");   -- @80 = 2 (compare_and_iter_f_init)

    -- Load signals for each cycle
      type t1load_data_array is array (natural range <>) of
         std_logic_vector(0 downto 0);

      constant t1load_data : t1load_data_array :=
      ("1",      -- @0 = 1
       "1",      -- @1 = 1
       "1",      -- @2 = 1
       "1",      -- @3 = 1
       "1",      -- @4 = 1
       "1",      -- @5 = 1
       "1",      -- @6 = 1
       "1",      -- @7 = 1
       "1",      -- @8 = 1
       "1",      -- @9 = 1
       "1",      -- @7 = 1
       "1",      -- @8 = 1
       "1",      -- @9 = 1
       "1",      -- @10 = 1
       "1",      -- @11 = 1
       "1",      -- @12 = 1
       "1",      -- @13 = 1
       "1",      -- @14 = 1
       "1",      -- @15 = 1
       "1",      -- @16 = 1
       "1",      -- @17 = 1
       "1",      -- @18 = 1
       "1",      -- @19 = 1
       "1",      -- @20 = 1
       "1",      -- @21 = 1
       "1",      -- @22 = 1
       "1",      -- @23 = 1
       "1",      -- @24 = 1
       "1",      -- @25 = 1
       "1",      -- @26 = 1
       "1",      -- @27 = 1
       "1",      -- @28 = 1
       "1",      -- @29 = 1
       "1",      -- @30 = 1
       "1",      -- @31 = 1
       "1",      -- @32 = 1
       "1",      -- @33 = 1
       "1",      -- @34 = 1
       "1",      -- @35 = 1
       "1",      -- @36 = 1
       "1",      -- @37 = 1
       "1",      -- @38 = 1
       "1",      -- @39 = 1
       "1",      -- @40 = 1
       "1",      -- @41 = 1
       "1",      -- @42 = 1
       "1",      -- @43 = 1
       "1",      -- @44 = 1
       "1",      -- @45 = 1
       "1",      -- @46 = 1
       "1",      -- @47 = 1
       "1",      -- @48 = 1
       "1",      -- @49 = 1
       "1",      -- @50 = 1
       "1",      -- @51 = 1
       "1",      -- @52 = 1
       "1",      -- @53 = 1
       "1",      -- @54 = 1
       "1",      -- @55 = 1
       "1",      -- @56 = 1
       "1",      -- @57 = 1
       "1",      -- @58 = 1
       "1",      -- @59 = 1
       "1",      -- @60 = 1
       "1",      -- @61 = 1
       "1",      -- @62 = 1
       "1",      -- @63 = 1
       "1",      -- @64 = 1
       "1",      -- @65 = 1
       "1",      -- @66 = 1
       "1",      -- @67 = 1
       "1",      -- @68 = 1
       "1",      -- @69 = 1
       "1",      -- @70 = 1
       "1",      -- @71 = 1
       "1",      -- @72 = 1
       "1",      -- @73 = 1
       "1",      -- @74 = 1
       "1",      -- @75 = 1
       "1",      -- @76 = 1
       "1",      -- @77 = 1
       "1",      -- @78 = 1
       "1",      -- @79 = 1
       "0");     -- @80 = 0

      type t2load_data_array is array (natural range <>) of
         std_logic_vector(0 downto 0);

      constant t2load_data : t2load_data_array :=
      ("1",      -- @0 = 1
       "1",      -- @1 = 1
       "1",      -- @2 = 1
       "1",      -- @3 = 1
       "1",      -- @4 = 1
       "1",      -- @5 = 1
       "1",      -- @6 = 1
       "1",      -- @7 = 1
       "1",      -- @8 = 1
       "1",      -- @9 = 1
       "1",      -- @7 = 1
       "1",      -- @8 = 1
       "1",      -- @9 = 1
       "1",      -- @10 = 1
       "1",      -- @11 = 1
       "1",      -- @12 = 1
       "1",      -- @13 = 1
       "1",      -- @14 = 1
       "1",      -- @15 = 1
       "1",      -- @16 = 1
       "1",      -- @17 = 1
       "1",      -- @18 = 1
       "1",      -- @19 = 1
       "1",      -- @20 = 1
       "1",      -- @21 = 1
       "1",      -- @22 = 1
       "1",      -- @23 = 1
       "1",      -- @24 = 1
       "1",      -- @25 = 1
       "1",      -- @26 = 1
       "1",      -- @27 = 1
       "1",      -- @28 = 1
       "1",      -- @29 = 1
       "1",      -- @30 = 1
       "1",      -- @31 = 1
       "1",      -- @32 = 1
       "1",      -- @33 = 1
       "1",      -- @34 = 1
       "1",      -- @35 = 1
       "1",      -- @36 = 1
       "1",      -- @37 = 1
       "1",      -- @38 = 1
       "1",      -- @39 = 1
       "1",      -- @40 = 1
       "1",      -- @41 = 1
       "1",      -- @42 = 1
       "1",      -- @43 = 1
       "1",      -- @44 = 1
       "1",      -- @45 = 1
       "1",      -- @46 = 1
       "1",      -- @47 = 1
       "1",      -- @48 = 1
       "1",      -- @49 = 1
       "1",      -- @50 = 1
       "1",      -- @51 = 1
       "1",      -- @52 = 1
       "1",      -- @53 = 1
       "1",      -- @54 = 1
       "1",      -- @55 = 1
       "1",      -- @56 = 1
       "1",      -- @57 = 1
       "1",      -- @58 = 1
       "1",      -- @59 = 1
       "1",      -- @60 = 1
       "1",      -- @61 = 1
       "1",      -- @62 = 1
       "1",      -- @63 = 1
       "1",      -- @64 = 1
       "1",      -- @65 = 1
       "1",      -- @66 = 1
       "1",      -- @67 = 1
       "1",      -- @68 = 1
       "1",      -- @69 = 1
       "1",      -- @70 = 1
       "1",      -- @71 = 1
       "1",      -- @72 = 1
       "1",      -- @73 = 1
       "1",      -- @74 = 1
       "1",      -- @75 = 1
       "1",      -- @76 = 1
       "1",      -- @77 = 1
       "1",      -- @78 = 1
       "1",      -- @79 = 1
       "0");     -- @80 = 0


    -- Arrays for expected outputs for each output port.
      type r1data_data_array is array (natural range <>) of
         std_logic_vector(31 downto 0);

      constant r1data_data : r1data_data_array :=
      ("00000000000000000000000000000000",       -- @0 = 0
       "00000000000000000010000000010000",       -- @1 = 8208 (compare_and_iter_f)
       "00000000000000000100100000011000",       -- @2 = 18456 (compare_and_iter_f)
       "00000000000000000010000011110000",       -- @3 = 8432 (compare_and_iter_f)
       "00000000001001110100101100010100",       -- @4 = 2575124  (compare_and_iter_f)
       "00000000001001110111111100011100",       -- @5 = 2588444 (compare_and_iter_f)
       "11111111110110010010101111101100",       -- @6 = -2544660 (compare_and_iter_f)
       "00000000001001111100001100100100",       -- @7 = 2605860 (compare_and_iter_f)
       "00000000000000000010000000010000",       -- @8 = 8208 (compare_and_iter_f)
       "00000000000000000100100000011000",       -- @9 = 18456 (compare_and_iter_f)
       "11111111110110001111101100001100",       -- @10 = -2557172  (compare_and_iter_f)
       "11111111110110010001011100010100",       -- @11 = -2549996 (compare_and_iter_f)
       "11111111110110010100001100011100",       -- @12 = -2538724    (compare_and_iter_f)
       "00000000001001110011011111101100",       -- @13 = 2570220 (compare_and_iter_f)



       "11010000100111011000110001011101",       -- @11 = 3499986013
       "11000100000111101010010110011110",       -- @12 = 3290342814
       "10111001011111110111101110110011",       -- @13 = 3112139699
       "11000011110100110110110001001101",       -- @14 = 3285412941
       "00101011101010011001110110000001",       -- @15 = 732536193
       "00010110001001001110001101000101",       -- @16 = 371516229
       "11001001010001011100101010001011",       -- @17 = 3376794251
       "10011001000000100101000111001001",       -- @18 = 2567066057
       "11100010101001111010100000000111",       -- @19 = 3802638343
       "01101101101110110011001000011011",       -- @20 = 1840984603
       "00010001110000000101111100111100",       -- @21 = 297819964
       "10011000010011000110100101101001",       -- @22 = 2555144553
       "10001101101011100100011100000000",       -- @23 = 2377008896
       "01101001101101111010011010000100",       -- @24 = 1773643396
       "01110000111100101011110101010110",       -- @25 = 1894956374
       "00011000000011001111100011000111",       -- @26 = 403503303
       "11010011110111100100110101010110",       -- @27 = 3554561366
       "01001001011010101001101110111111",       -- @28 = 1231723455
       "10000100000101100000010101100011",       -- @29 = 2216035683
       "11110111001011111011110101111110",       -- @30 = 4147101054
       "11110101011110101101111011010110",       -- @31 = 4118470358
       "01111101111110010100111110010001",       -- @32 = 2113490833
       "10101110001100010101110111110000",       -- @33 = 2922470896
       "00110001010100100100010110010010",       -- @34 = 827475346
       "10010000010001000010101001110011",       -- @35 = 2420386419
       "01000011001101001111111001010000",       -- @36 = 1127546448
       "01011111010101110000100100010100",       -- @37 = 1599539476
       "00111010001101001110010001111011",       -- @38 = 976544891
       "10101010001100110000000111101000",       -- @39 = 2855469544
       "10000011101000000100101110001000",       -- @40 = 2208320392
       "01101010000100011000110110100001",       -- @41 = 1779535265
       "10000001111110010010011110110110",       -- @42 = 2180589494
       "00110110001010000111001001100011",       -- @43 = 908620387
       "11110100010011110100101110001001",       -- @44 = 4098837385
       "10100000111100110100101100100010",       -- @45 = 2700299042
       "01001000111001111011110111101000",       -- @46 = 1223146984
       "01011101001111110001100000101011",       -- @47 = 1564416043
       "11000000000100101011011001011110",       -- @48 = 3222451806
       "11001101111100011000011110100000",       -- @49 = 3455158176
       "01110110111110001001001110111100",       -- @50 = 1996002236
       "11110101111000000010001101010010",       -- @51 = 4125107026
       "10010010100000111001100111100000",       -- @52 = 2458098144
       "01111101011101001101000010001101",       -- @53 = 2104807565
       "00011101000011010011101011111100",       -- @54 = 487406332
       "01010000010000001100110100010111",       -- @55 = 1346424087
       "10000000111100001111010101010000",       -- @56 = 2163275088
       "10001010001111110100111001011110",       -- @57 = 2319404638
       "11110000111101111000101100010110",       -- @58 = 4042754838
       "10110101111111010111111101110000",       -- @59 = 3053289328
       "11111110010100010000001010011111",       -- @60 = 4266721951
       "11101001011100010001011101000000",       -- @61 = 3916502848
       "10001110100011000101001011101001",       -- @62 = 2391560937
       "00010110010011000001101010001101",       -- @63 = 374086285
       "11100100111111011101111101010010",       -- @64 = 3841843026
       "11001001111111111111001110101011",       -- @65 = 3388994475
       "11110000010000001001010000100011",       -- @66 = 4030764067
       "00111011010001000001001110111111",       -- @67 = 994317247
       "10110110111000001100010111110001",       -- @68 = 3068184049
       "10000100101111110000010010101111",       -- @69 = 2227111087
       "11101010111101010000100001101110",       -- @70 = 3941927022
       "00000000000000000000000000000000",       -- @71 = 2213459199
       "00000000000000000001001000000100",       -- @72 = 1454268293
       "00000000000000000100011000010100",       -- @73 = 1614888088
       "11111111111111110111110000011000",       -- @74 = 2241593203
       "00000000000000011011100000101000",       -- @75 = 2740546453
       "11111111111111011110010001001000",       -- @76 = 4255533836
       "00000000000000100010000001000100",       -- @77 = 1870913602
       "11111111111111111100000000100000",       -- @78 = 3181588603
       "00000000000000101010110001001000",       -- @79 = 50739021
       "00000000000000010000111000111100"        -- @80 = 725711285
        );     

      constant IGNORE_OUTPUT_COUNT : integer := 1;
      constant TOTAL_CYCLE_COUNT : integer := 81;


     variable current_cycle : integer;
  begin

    -- Initialize the clock signal.
    clk <= '0';

    -- Reset active to initialize regs
    rstx <= '0';
    wait for 1 ns;

    -- Release reset.
    rstx <= '1';
    -- Global lock off.
    glock <= '0';


    for current_cycle in 0 to TOTAL_CYCLE_COUNT - 1 loop

    -- The actual test bench code.
      t1data <= t1data_data(current_cycle);
      t1load <= t1load_data(current_cycle);
      t2data <= t2data_data(current_cycle);
      t2load <= t2load_data(current_cycle);
      t1opcode <= t1opcode_data(current_cycle);

      if current_cycle >= IGNORE_OUTPUT_COUNT then
         assert r1data = r1data_data(current_cycle)
            report lf & "TCE Assert: Verification failed at cycle " & integer'image(current_cycle) & " for output 0"
            & " actual: " & integer'image(to_integer(signed(r1data)))
            & " expected: " & integer'image(to_integer(signed(r1data_data(current_cycle))))  severity error;

      end if;

      -- Generate a clock pulse.
      -- TODO: Generate the clock in a separate component.
      wait for 1 ns;
      clk <= not clk;
      wait for 1 ns;
      clk <= not clk;

    end loop;  -- current_cycle

    -- Ends the simulation (at least in case of ghdl).
    wait;
  end process;
end behav;